----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:37:56 12/05/2017 
-- Design Name: 
-- Module Name:    VGA_game_control - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity VGA_game_control is
                 port(
							clk_25m:in std_logic;
							rst_n:in std_logic;
							key_signal : in std_logic;--------�м�ֵ���µı�־λ
							ps2_data: in std_logic_vector(7 downto 0);
							is_moving:out std_logic_vector(8 downto 0);
							game_score:out std_logic_vector(7 downto 0)
	    
					      );
end VGA_game_control;

architecture Behavioral of VGA_game_control is
constant time_1s:integer:=24999999;
constant time_0p5s:integer:= 12499999;
constant time_0p25s:integer:= 6249999;
constant updata_coordinate_time:integer:=49999;
signal fresh_time:integer range 0 to 50000000:=24999999;
signal fresh_time_cnt:integer range 0 to 50000000:=0;
signal game_score_temp:std_logic_vector(7 downto 0);
signal is_moving_temp:std_logic_vector(8 downto 0);
signal body_cnt:integer range 0 to 8:=0;
signal body_set1:integer range 0 to 8:=0;
signal body_set2:integer range 0 to 8:=0;
signal m_sequence:std_logic_Vector(5 downto 0):="11"&X"F";
signal updata_time:integer range 0 to 24999999:=0;
begin
game_score<=game_score_temp;
is_moving<=is_moving_temp;
refresh_pro:process(clk_25m,rst_n)
begin
    if rst_n='0' then
	  fresh_time<=time_1s;
	elsif rising_edge(clk_25m)then
       if game_score_temp<=X"09" then
		   fresh_time<=time_1s;
	    elsif game_score_temp>X"09" and game_score_temp<=	X"19" then
		   fresh_time<=time_0p5s;
		 elsif game_score_temp>X"19" then
		   fresh_time<=time_0p25s;
		end if;
	end if;	
end  process refresh_pro;


score_ctrl:process(clk_25m,rst_n)
begin
   if rst_n='0' then
	   game_score_temp<=X"00"; 
	elsif	rising_edge(clk_25m) then
	   if key_signal='1' and is_moving_temp(conv_integer(ps2_data(3 downto 0)))='1' then
            if game_score_temp(3 downto 0)=X"9" then
				    if game_score_temp(7 downto 4)=X"9" then
					      game_score_temp<=X"00";
					 else
				         game_score_temp(7 downto 4)<=game_score_temp(7 downto 4)+1;
					     	game_score_temp(3 downto 0)<=X"0";
					 end if;		
				else
				  game_score_temp(3 downto 0)<=game_score_temp(3 downto 0)+1;
				end if; 
   end if;
end if;	
end process score_ctrl;



body_cnt_ctrl:process(clk_25m,rst_n)
begin
    if rst_n ='0' then
	    body_cnt<=0;
	 elsif rising_edge(clk_25m) then
       if body_cnt=8 then
	  	   body_cnt<=0;
		 else
		   body_cnt<=body_cnt+1;
		end if;
	end if;	
end process body_cnt_ctrl;

process(clk_25m,rst_n)
begin
    if rst_n='0' then
	    fresh_time_cnt<=0;
	 elsif rising_edge(clk_25m)	then
      if fresh_time_cnt>=fresh_time then
        	fresh_time_cnt<=0;
		else
	      fresh_time_cnt<=fresh_time_cnt+1;
		end if;
end if;		
end process;


process(clk_25m,rst_n)
begin
   if rst_n='0' then
	     is_moving_temp<=(others=>'0');
	elsif rising_edge(clk_25m)	then
    	if fresh_time_cnt=fresh_time and  game_score_temp<=X"09" then
		   case(body_set1) is
			    when 0=>
				         is_moving_temp(0)<='1';
							is_moving_temp(7 downto 1)<=(others=>'0');
		       when 1=>
				         is_moving_temp<=(1=>'1',others=>'0');
			    when 2=>
				         is_moving_temp<=(2=>'1',others=>'0');	
			    when 3=>
				         is_moving_temp<=(3=>'1',others=>'0');
			    when 4=>
				         is_moving_temp<=(4=>'1',others=>'0');	
			    when 5=>
				         is_moving_temp<=(5=>'1',others=>'0');	
			    when 6=>
				         is_moving_temp<=(6=>'1',others=>'0');	
			    when 7=>
				         is_moving_temp<=(7=>'1',others=>'0');	
             when others=>null;
			end case;	 
      elsif	fresh_time_cnt=fresh_time and  game_score_temp>X"09" then
          case(body_set1) is
			    when 0=>
						   is_moving_temp<=(1=>'1',7=>'1',others=>'0');
		       when 1=>
				         is_moving_temp<=(1=>'1',3=>'1',others=>'0');
			    when 2=>
				         is_moving_temp<=(2=>'1',1=>'1',others=>'0');	
			    when 3=>
				         is_moving_temp<=(3=>'1',5=>'1',others=>'0');
			    when 4=>
				         is_moving_temp<=(4=>'1',7=>'1',others=>'0');	
			    when 5=>
				         is_moving_temp<=(5=>'1',2=>'1',others=>'0');	
			    when 6=>
				         is_moving_temp<=(6=>'1',8=>'1',others=>'0');	
			    when 7=>
				         is_moving_temp<=(7=>'1',4=>'1',others=>'0');	
             when others=>null;
			end case;	      		
		  else
        is_moving_temp<=is_moving_temp;
	   end if;
end if;		
end process;


process(clk_25m,rst_n)
begin
   if rst_n='0' then
	  m_sequence<="11"&X"F";
	elsif rising_edge(clk_25m)	then
	  m_sequence<=(m_sequence(0) xor m_sequence(1))&m_sequence( 5 downto 1);
	end if;  
end process;


process(clk_25m,rst_n)
begin
   if rst_n='0' then
	   updata_time<=updata_coordinate_time;
	elsif rising_edge(clk_25m)	then
       if fresh_time_cnt=fresh_time  then
	  	 updata_time<=updata_coordinate_time+conv_integer(m_sequence);
		 else
		 updata_time<=updata_time;
		 end if;
end if;		 
end process;



process(clk_25m,rst_n)
begin
   if rst_n='0' then
	   body_set1<=0;
   elsif rising_edge(clk_25m)	then
   if fresh_time_cnt=updata_time then
      body_set1<=body_cnt;
    else
      body_set1<=body_set1;
  end if;
end if;  
end process;
end Behavioral;

